/*
Write a markdown documentation for this systemverilog module:
Author : S. M. Tahmeed Reza (https://github.com/tahmeedKENJI)
This file is part of DSInnovators:rv64g-core
Copyright (c) 2024 DSInnovators
Licensed under the MIT License
See LICENSE file in the project root for full license information
*/

module pipeline_lite #(
    parameter int DATAWIDTH = 32
) (
    input logic arst_ni,
    input logic clk_i,
    input logic clear_i,
    input logic [DATAWIDTH-1:0] data_in_i,
    input logic data_in_valid_i,
    output logic data_in_ready_o,
    output logic [DATAWIDTH-1:0] data_out_o,
    output logic data_out_valid_o,
    input logic data_out_ready_i
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS GENERATED
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  logic buffer_clear_flag;
  logic [DATAWIDTH-1:0] data_buffer;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  assign data_in_ready_o  = arst_ni & ~clear_i & ((buffer_clear_flag) ? '1 : data_out_ready_i);
  assign data_out_valid_o = arst_ni & ~clear_i & ~buffer_clear_flag;


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  always_ff @(posedge clk_i) begin
    if (~arst_ni) begin
      buffer_clear_flag <= '1;
    end else begin

      if (data_out_valid_o & data_out_ready_i) begin
        data_out_o <= data_buffer;
        buffer_clear_flag <= '1;
      end
      if (data_in_valid_i & data_in_ready_o) begin
        data_buffer <= data_in_i;
        buffer_clear_flag <= '0;
      end

    end
  end

  // always_ff @( posedge clk_i or negedge arst_ni ) begin : blockName
  //   if (data_in_ready_o & data_in_valid_i) begin
  //     data_out_o <= data_in_i;
  //   end
  // end
  // always_ff @(posedge clk_i) begin
  //   if (~arst_ni) buffer_clear_flag <= '1;
  //   else begin
  //     casex ({
  //       clear_i, data_in_valid_i, data_in_ready_o, data_out_valid_o, data_out_ready_i
  //     })
  //       5'b1xxxx, 5'b00011: buffer_clear_flag <= '1;
  //       5'b01100, 5'b01111: buffer_clear_flag <= '0;
  //       default: buffer_clear_flag <= buffer_clear_flag;
  //     endcase
  //   end
  // end

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INITIAL CHECKS
  //////////////////////////////////////////////////////////////////////////////////////////////////

`ifdef SIMULATION
  initial begin
    if (DATAWIDTH > 2) begin
      $display("\033[1;33m%m DATAWIDTH\033[0m");
    end
  end
`endif  // SIMULATION

endmodule
